`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:10:28 09/11/2022 
// Design Name: 
// Module Name:    adder_carry_95_Amisha 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder_carry_95_Amisha(a_amisha, b_amisha, sum_amisha, cout_amisha);
	 parameter N = 4;
	 parameter N1 = N-1;
    input wire [N1:0] a_amisha;
    input wire [N1:0] b_amisha;
    output wire [N1:0] sum_amisha;
    output cout_amisha;
	 
	 wire [N:0] sum_ext_amisha;
	 
	 assign sum_ext_amisha = {1'b0, a_amisha} + {1'b0, b_amisha};
	 assign sum_amisha = sum_ext_amisha[N1:0];
	 assign cout_amisha = sum_ext_amisha[N];
endmodule
